module decoder_3_to_8_1202212ferdous (
input [2:0] C,
output [7:0] O
);
assign O = (C == 3'b000) ? 8'b00010001 :
(C == 3'b001) ? 8'b00100010 :
(C == 3'b010) ? 8'b01000100 :
(C == 3'b011) ? 8'b10000100 :
(C == 3'b100) ? 8'b00010000 :
(C == 3'b101) ? 8'b00001000 :
(C == 3'b110) ? 8'b00000100 :
8'b00000010;
endmodule
